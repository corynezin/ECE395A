with adr select sel <=
	d(0) when "0000000",
	d(1) when "0000001",
	d(2) when "0000010",
	d(3) when "0000011",
	d(4) when "0000100",
	d(5) when "0000101",
	d(6) when "0000110",
	d(7) when "0000111",
	d(8) when "0001000",
	d(9) when "0001001",
	d(10) when "0001010",
	d(11) when "0001011",
	d(12) when "0001100",
	d(13) when "0001101",
	d(14) when "0001110",
	d(15) when "0001111",
	d(16) when "0010000",
	d(17) when "0010001",
	d(18) when "0010010",
	d(19) when "0010011",
	d(20) when "0010100",
	d(21) when "0010101",
	d(22) when "0010110",
	d(23) when "0010111",
	d(24) when "0011000",
	d(25) when "0011001",
	d(26) when "0011010",
	d(27) when "0011011",
	d(28) when "0011100",
	d(29) when "0011101",
	d(30) when "0011110",
	d(31) when "0011111",
	d(32) when "0100000",
	d(33) when "0100001",
	d(34) when "0100010",
	d(35) when "0100011",
	d(36) when "0100100",
	d(37) when "0100101",
	d(38) when "0100110",
	d(39) when "0100111",
	d(40) when "0101000",
	d(41) when "0101001",
	d(42) when "0101010",
	d(43) when "0101011",
	d(44) when "0101100",
	d(45) when "0101101",
	d(46) when "0101110",
	d(47) when "0101111",
	d(48) when "0110000",
	d(49) when "0110001",
	d(50) when "0110010",
	d(51) when "0110011",
	d(52) when "0110100",
	d(53) when "0110101",
	d(54) when "0110110",
	d(55) when "0110111",
	d(56) when "0111000",
	d(57) when "0111001",
	d(58) when "0111010",
	d(59) when "0111011",
	d(60) when "0111100",
	d(61) when "0111101",
	d(62) when "0111110",
	d(63) when "0111111",
	d(64) when "1000000",
	d(65) when "1000001",
	d(66) when "1000010",
	d(67) when "1000011",
	d(68) when "1000100",
	d(69) when "1000101",
	d(70) when "1000110",
	d(71) when "1000111",
	d(72) when "1001000",
	d(73) when "1001001",
	d(74) when "1001010",
	d(75) when "1001011",
	d(76) when "1001100",
	d(77) when "1001101",
	d(78) when "1001110",
	d(79) when "1001111",
	d(80) when "1010000",
	d(81) when "1010001",
	d(82) when "1010010",
	d(83) when "1010011",
	d(84) when "1010100",
	d(85) when "1010101",
	d(86) when "1010110",
	d(87) when "1010111",
	d(88) when "1011000",
	d(89) when "1011001",
	d(90) when "1011010",
	d(91) when "1011011",
	d(92) when "1011100",
	d(93) when "1011101",
	d(94) when "1011110",
	d(95) when "1011111",
	d(96) when "1100000",
	d(97) when "1100001",
	d(98) when "1100010",
	d(99) when "1100011",
	d(100) when "1100100",
	d(101) when "1100101",
	d(102) when "1100110",
	d(103) when "1100111",
	d(104) when "1101000",
	d(105) when "1101001",
	d(106) when "1101010",
	d(107) when "1101011",
	d(108) when "1101100",
	d(109) when "1101101",
	d(110) when "1101110",
	d(111) when "1101111",
	d(112) when "1110000",
	d(113) when "1110001",
	d(114) when "1110010",
	d(115) when "1110011",
	d(116) when "1110100",
	d(117) when "1110101",
	d(118) when "1110110",
	d(119) when "1110111",
	d(120) when "1111000",
	d(121) when "1111001",
	d(122) when "1111010",
	d(123) when "1111011",
	d(124) when "1111100",
	d(125) when "1111101",
	d(126) when "1111110",
	d(127) when "1111111";
