PACKAGE data_types is
	
	type conv_0_input is array (0 to 2) of signed(7 downto 0);
	type conv_0_output is array (0 to 3) of signed (7 downto 0);

END data_types;
