
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package arrays is
type output_array is array (0 to 63) of STD_LOGIC_VECTOR(47 downto 0);
end arrays;