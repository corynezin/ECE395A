package body MATRIX is
constant matrix_height: INTEGER:= 100;
constant matrix_width: INTEGER:= 784;
constant number_size: INTEGER:= 8;
end MATRIX;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use WORK.MATRIX.ALL;
package vector_v is
constant v: vector_in:=(
"11100000","01010110","11100000","01010000","00100000","01111101","10011111","00101011","10101110","11110110","10000111","10101000","10001011","11001101","00011010","10110110","10000111","00011100","01000000","11101010","10001000","11111101","00110001","00100001","00001011","01101001","11110011","00110010","10100001","01110111","11101100","01011011","00100110","11101100","00010100","00010011","11001110","11011000","11011000","00110100","00011110","00100010","11110100","11111001","11100110","10101000","10010010","00011011","10001111","10100111","11001000","10101001","01000010","00010011","00110110","10110101","11101000","10100100","01011100","10110111","11101010","10011101","01111110","01000100","11000100","00001001","11101101","00110111","11011100","01000010","01100100","10010101","00010010","00110011","11111101","01110000","00100011","00110110","10101101","10000000","00111001","10001111","01110011","10111000","00000010","01100101","00000011","01100111","10011101","00011010","10010101","00101010","01011111","10011011","01010100","00010000","00110010","11010101","10111000","00101100","01011101","11111000","01010111","00010100","11101101","00111100","10111001","01011101","00111111","10001101","00000101","11111010","00100011","11000011","10010100","01000111","01110001","10100001","11011101","10111101","01001000","10001010","01101100","01101000","10100110","10111000","00010110","01101001","00001110","01000100","10000101","11111110","01001010","01111000","00110011","01101100","01010001","01101101","00110001","11010000","10001100","01100101","00000010","01100101","00101011","10100010","10101111","10100101","00000010","11010010","01011100","01110111","01011000","00111011","10010111","00101101","00001010","00011011","10101010","01101001","00011010","11111110","00011001","00101100","11011010","00101100","10010010","01001011","11100111","11111110","11101010","01111101","00001100","00000010","10010100","01101101","11100000","11110000","10000101","11010111","11011110","11101101","11100110","01001111","00001100","11111110","10101001","11110101","10010010","10001000","01101011","00001001","01110000","00111110","01111100","10010111","11000111","10001000","11111110","11100010","00000001","11010101","00110010","00111001","11111100","10111011","11010010","00001011","11010000","10000100","00111110","11010100","10000001","01001100","00110011","00101000","00111011","00110011","01001001","11011100","11001110","00110100","11100010","11110111","10000100","01010000","00110011","00100001","10011010","01001011","01001110","11001111","00000100","10100111","00101111","10010110","10110100","10101001","10100011","01010111","00111100","00000100","01101100","00100111","01111000","11110101","01001111","01010101","01100100","11000011","11101011","00101000","10011000","00010100","11001101","11111101","00010111","00011101","00010101","10101000","01010101","10110110","01110101","01100110","10000100","00110110","00011001","00111101","10111101","11000001","01010100","00001010","01111101","00011001","10100000","11010011","11011101","01011000","00111111","11011100","00010101","10011010","00010100","11001011","00111010","11001110","01100011","01000010","00100011","01110111","11100110","11001010","11101111","11110100","01010001","11010111","01000101","01100101","01001100","10000110","10001111","00010011","10000110","10010001","10100100","01000011","00010111","10000111","00110011","01110110","01110001","10110110","00100111","11110000","10000010","01000001","00011100","11010110","00001011","01100111","00001101","10000100","01011111","00101011","01110110","01001000","11011010","01001010","11000110","01111010","10000000","10010101","11111000","11000011","00110001","11010001","00111001","11000100","10000100","01011111","10111101","11111100","10011110","01010110","01011011","11011001","00001001","11000101","10111000","01011110","00101100","01101010","11111111","10111000","11111011","01111000","01001000","11111010","01010000","11010110","10110001","11111001","11101010","00111110","11000011","10010100","00011001","01010101","11001001","11101111","01110011","00011101","11111101","10010111","11110011","00101101","00001010","11110101","00000100","00000001","10111100","11101000","10111000","10100011","11001110","11101111","01001001","10111000","11000100","10011010","01100111","11011111","01101000","11000001","11100100","10001110","10100111","00000101","01111011","00010011","10010100","01010010","10000100","01001110","01100110","00111110","10111111","00000001","01010011","00011101","11100110","01010001","01001000","11010110","11001111","01000001","00100000","10101111","11001101","00110100","10100010","10000101","11110010","00001101","11010101","01101100","00101110","10111001","11011010","10011011","01001010","00000100","11111000","01001000","01001000","01110110","00100010","10001101","10100111","11001000","01011110","00110000","01100111","11010110","00101101","11110101","11011111","00111101","11000110","11100110","00110000","00010010","00000001","11100011","10010010","11100010","11001101","01000110","01001101","11010000","10000011","10010110","11011101","11010001","11000111","00000011","01110111","10010110","11011000","00111010","10010100","00000100","10011110","00111100","00110111","00001010","00111101","00010111","11010001","11010110","10101111","10011001","00100100","11010101","00010110","10011011","10000100","00011100","00110111","10000011","11101101","11001111","00001101","01000001","00011110","01001110","00110101","11000100","01100110","01010100","11001101","10111101","10110010","10000010","01011111","10000100","01001110","01100000","00101000","00110101","10011100","00100110","10110111","00101100","01111101","00110100","11011000","01001011","01111101","11011010","10101110","11101001","00100110","10111000","00101000","10101011","01000110","11111100","10100001","01110101","10001100","00101101","10001100","01000100","10000010","10011110","00010001","00010011","11010100","11110110","01100111","10001011","11111101","00010000","11111100","01101100","01001010","00001111","01001010","10110010","11011110","10111110","00101001","11011001","00011001","00010100","01000111","10010101","00100001","10100000","01110011","11001000","01010011","00001010","10000100","01000000","11010101","11011000","00111000","00011111","11000001","00010010","10101101","00100011","10111011","01111101","01010011","11110111","11010100","01001000","01110101","11011000","11010100","11010100","11101100","11110010","10111001","00101011","01101010","11100000","01101100","11110001","11110111","00010010","10111001","10110011","11011110","00010110","10000111","01000111","10011011","10010101","01100010","11111111","10110111","11000100","01011001","01001110","01100010","00010111","01110111","10101101","00101110","10100111","11010001","01110100","11111011","01111010","01001010","10011101","11100001","11010101","11100000","11100011","10000110","11010000","00101011","10011000","10111110","11011010","01100110","11010010","10101010","01100011","11101111","11111001","01110000","01000011","01011000","11101110","00111000","01111100","11111100","10111001","10101000","00100111","01111110","00001101","01000111","00000111","01111110","11101111","10011101","10110110","10100011","01010101","10110000","10111101","11111011","10010101","11011010","00011001","01000110","10001100","10101011","01101011","10110001","01111101","01011000","11100100","00001001","01100011","01110011","01001100","00110010","10111000","00101101","10010110","10110111","01101100","10110101","10001000","01011101","00110100","10101111","11110011","10010011","00001000","00110011","00111011","11000111","01110110","01111100","01011000","10101001","11101001","11100011","11111011","11001111","01100101","10101010","01101110","11000110","11001001","00111001","10101110","00111111","11111010","10101110","01000110","10101011","11011001","01011000","11000001","10110110","01110110","00111010","10010010","01000100","00001100","11001100","00100001","10110111","11111101","10000101","00011111","00111100","00011010","00101101","00101011","11000101","01000001","11001010","10001110","11010110","00101011","10100100","00100001","01110111","11100000","00100001","00101111","01111110","00110110","11101111","11000000","11001001","01100101","11001011","01010100","11111111","10110101","01000011","11000010","10100001","00100001","01011110","11001100","11011001","00101011","11101001","01001010","00010100","00111111","10000110","00100101","10111010","01100011","10010010","01010011","01110110","10011001","11100010","01111100","11011111","11101111","10101000","00101010","01101001","11100001","01111011","11001010","01011001","11111000");
end package;