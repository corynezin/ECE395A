package body MATRIX is
constant matrix_height: INTEGER:= 100;
constant matrix_width: INTEGER:= 784;
constant number_size: INTEGER:= 8;
end MATRIX;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use WORK.MATRIX.ALL;
package vector_w is
constant w: vector_in:=(
"00000010","01000110","11001001","01110001","00000011","11110010","01101011","10101000","11010101","00010001","01101101","11010100","11100110","01001011","01000111","10010101","10110111","11111101","01110100","11011010","01110111","00110000","01110110","00001000","10010110","10110100","10000111","10100001","11001000","00101010","00000011","10001001","00001011","01000111","00100111","11011101","00111111","10000100","11101010","01000100","01101000","10010101","10110111","10001100","00001000","11111111","11111011","01101011","00001011","11110101","10011111","01110001","01011000","10100011","01001100","01001010","11111000","00111011","11101100","10011100","01011000","10100111","00010011","00011011","01110100","10100100","10010100","10100100","10101100","10010100","11111001","11100100","11111101","10000000","00100100","10001001","11010001","11100001","01011101","10010111","00011101","01000110","11000101","11000001","01001000","00011100","01011001","01110010","00000110","01101001","00011100","01001011","11101101","11001001","01110101","11100001","00001000","10111100","11001000","01110010","10010100","01100000","01000010","11110110","00010000","00100010","11101101","00111101","01011101","00000000","00011000","11010110","10111010","10100111","01101001","11010110","00101000","00010100","11110111","00010111","01110110","10100101","11010100","11100111","10110100","11100000","10101001","11001111","10110010","11001101","01001000","11001001","11111101","01111101","00101101","10011011","11111001","01011000","10110011","10000100","11111111","00000100","00100000","10010101","10111001","01001110","00010100","00110010","00000101","11000011","11000010","11100001","11010111","00111011","11001101","11001011","10110011","01000101","00011010","11110011","11010001","01001110","11011100","01111010","00010111","01001010","00010100","00111011","11000000","11100001","10000011","01111101","01011111","01101011","00111100","01101001","00111100","00101010","11010011","00001011","01010100","01010001","11010110","10011101","00100101","10110010","11000000","01001101","10010010","11111110","11001101","10001111","11010010","00111100","00100101","10101100","10111100","10101010","01101011","11001001","11101111","11010011","10101010","10010100","00011011","00100111","11011110","10011110","00100110","11111111","10111011","11010110","11100100","00001000","00001011","00111111","11101101","10100111","00001111","11011001","01101101","11100100","11100101","01010111","10000100","11100011","10000111","10010000","10011110","11001010","00111000","00011001","00111110","11000100","10101111","11000010","00000010","01010100","10010010","01000000","00111011","00101101","10010011","10101010","10010100","00000111","10010101","10110000","00010010","10000011","01011011","11110010","11100000","10011001","10001111","10110010","00110011","00001110","11111010","01011000","00101010","11100101","01101011","01011000","00011011","00111010","00001110","10001101","00101000","01001110","10110000","10000100","10111010","01110011","01101000","01000101","01111011","01111101","01000000","11110010","10001111","01110110","00111010","11000000","11110110","00011110","11110000","11101001","01010100","01000111","11000100","11010001","00001001","10001010","01010101","01100100","00001000","00011001","10000101","11011101","11101011","00110011","00011111","11100101","01011101","10001111","11010000","11111111","01011011","10000011","10000010","00110011","01100100","00110001","01011010","11000100","10110011","10010010","00111110","10010001","00101111","01110100","01100100","11011101","01001110","00100010","00111101","01011111","10010110","00000111","01001011","11010110","01000011","11000101","01101001","11110011","10101110","11010001","00001011","10001010","11110011","10001001","10110011","10111010","11100100","00011011","11010011","10100011","00100001","11111100","00100111","00010010","10111011","01010010","01001101","00111100","11011111","11000101","10001010","11101001","00101000","01001100","10110110","00110101","11001111","11100001","00100101","11101101","11110000","01000001","11111011","11111010","01010000","00000101","11001111","01100110","10101100","11110100","10010000","00110100","11000100","11111110","11101110","00101111","01111101","11110100","00111100","00010011","10011100","11110101","01110011","00010100","00011001","10011110","10110001","00111101","11110000","11011101","11001111","10111111","10101010","01111000","01100001","01110110","01001001","10110000","10000000","10011000","10100100","00110101","01101101","10001101","10000101","00000110","11011110","01011010","10101110","00110000","10001000","11000010","11110001","00011111","11010001","11000000","10001010","01001111","00110000","01100011","11001000","01111001","10010001","11111101","11110011","11110010","11110010","10111010","01111011","00000110","00100111","00110111","01100110","01100011","11010011","11011001","10010110","11100011","10101110","00001101","00100100","10011011","00100110","11110111","11100000","11001011","10011110","10110011","11110111","01010000","01101110","10000110","01010100","00011101","11110001","00010100","11011101","10101011","01110010","01111010","01110001","01100000","10101001","11011100","01001111","11101111","00011110","10110110","10110111","11001101","10000000","01001101","01100011","11101101","01010111","01011101","01101101","01000011","00010010","01010001","01110111","01110101","01111111","10110101","11001100","10111001","11010101","00011000","01110000","00010011","01101111","01100011","00110100","11110000","11101000","01100101","00111010","10111000","01000011","00111101","10001100","01010000","10101111","01100010","10100111","10011000","01111010","00010100","01110010","10110010","10100001","01101111","00101001","11111100","01110000","00111110","01000101","11001001","11010111","00010000","10010101","10001101","11110011","11110011","11111101","11100111","01010000","10001100","11101011","11100011","01000000","11100000","10001111","11111000","00101000","01001110","01101010","00111110","11011100","11101101","01001011","01100101","01001010","10010001","10000011","11101111","00110011","00010001","10110111","10111101","00110010","10100001","10111110","00100000","01001011","10011001","11100101","11010011","01111101","01101101","01010111","01110001","01011000","10110001","10000111","00000100","11110100","10010011","11011000","11111111","00011010","10100110","11100100","00010000","00100101","10110101","11110100","10001100","11100011","10101110","11011011","01111100","10111101","00000100","10100000","01110100","00010111","11001111","10000111","00101100","01110110","01101000","00001010","00000001","01010111","01111001","01011111","10101100","11000000","11101111","01100011","00001011","11000101","01101110","01100001","00010001","11010001","10100001","01010111","10110101","00100011","10000011","01000011","01000010","01110101","00111011","01100101","01111100","10000001","11100001","00100100","00011100","01001100","10001000","00000011","10101011","00000111","10000110","10110000","10100000","11000101","00000101","11111001","10100001","11010101","00100001","10010010","01000100","10111100","00010010","10011101","10110011","01110110","10011010","01110111","11011010","01101100","11100101","01111010","00110111","01010110","11110000","00010010","11011011","10000100","10001111","01001100","10001010","00101010","11100111","00010100","00001011","00001001","11101100","00101001","00111011","01100001","00101101","01000010","00001011","00001011","01001001","11110011","10000110","00101101","11111000","11011100","00001100","10011110","01111001","01100011","01001100","10101010","01011101","00010000","01011110","00010000","11000101","00000010","11011111","10001010","01010100","00010100","10110111","00110110","00010011","11101010","00111010","01011001","10001010","10100111","11110111","10100010","11111000","11111100","10010111","00001101","11101001","11000010","11010010","01011100","00110001","11110111","11110111","00101101","10001110","11000010","00100010","11000101","00011011","11110111","11010001","11011011","10101010","00110001","11011101","01000101","00111101","11001111","10111001","00010110","00010100","11101101","01111111","01111110","01011100","11001000","00101101","00100010","10011110","10110101","00100010","11110110","10110110","10010110","10101110","11001000","01110010","00101100","11101001","00011101","01101011","00111110","11100110","00110111","11100001","00100010","01110110","10010101","11110000","11111101","01001000","00111001","11000001","00110111","10010011","10100011","00101001","01110111","10101001","01101010","11001111","00111010","11111110","00000110","00111101");
end package;